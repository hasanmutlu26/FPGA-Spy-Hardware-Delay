// Causes direct delay. 

module singlepath_3 (N11334, N251);
(* keep = 1 *) input N251;
(* keep = 1 *) output N11334;
(* keep = 1 *) wire N11313, N11278, N11260, N11321, N11213, N11168, N11115, N11299, N11044, N10988, N10872, N10737, N11328, N10671, N5683, N10672, N6779, N9067, N4471, N1990, N1302, N11242, N3114, N3515, N6783, N9957, N3149, N10989, N10928, N644, N10873, N643, N11314, N6773, N7465, N11114, N6762, N10314, N1833, N8114, N10789, N10509, N10170, N9432, N9066, N10315, N9642, N11214, N9958, N1323, N5171, N7447, N10431;


buf BUFF1_58(N643, N251);
not NOT1_59(N644, N251);
buf BUFF1_162(N1302, N644);
buf BUFF1_169(N1323, N644);
not NOT1_262(N1833, N1302);
and AND2_351(N1990, N644, 1'b1);
and AND2_680(N3114, N644, 1'b1);
and AND2_691(N3149, N644, 1'b1);
nor NOR2_786(N3515, N644, 1'b0);
nand NAND2_939(N4471, N1833, 1'b1);
nand NAND2_1282(N5171, N1302, 1'b1);
nand NAND2_1394(N5683, N4471, 1'b1);
and AND5_1750(N6762, N5683, 1'b1, 1'b1, 1'b1, 1'b1);
and AND4_1758(N6773, N5683, 1'b1, 1'b1, 1'b1);
and AND3_1764(N6779, N5683, 1'b1, 1'b1);
and AND2_1768(N6783, N5683, 1'b1);
buf BUFF1_1959(N7447, N5683);
buf BUFF1_1965(N7465, N5683);
or OR4_2030(N8114, N6779, 1'b0, 1'b0, 1'b0);
not NOT1_2398(N9066, N8114);
nand NAND2_2399(N9067, N8114, 1'b1);
nand NAND2_2552(N9432, N9066, 1'b1);
nand NAND2_2648(N9642, N9432, 1'b1);
not NOT1_2793(N9957, N9642);
nand NAND2_2794(N9958, N9642, 1'b1);
nand NAND2_2919(N10170, N9958, 1'b1);
not NOT1_2987(N10314, N10170);
nand NAND2_2988(N10315, N10170, 1'b1);
nand NAND2_3032(N10431, N10314, 1'b1);
nand NAND2_3049(N10509, N10431, 1'b1);
not NOT1_3138(N10671, N10509);
nand NAND2_3139(N10672, N10509, 1'b1);
nand NAND2_3181(N10737, N10671, 1'b1);
nand NAND2_3212(N10789, N10737, 1'b1);
not NOT1_3254(N10872, N10789);
nand NAND2_3255(N10873, N10789, 1'b1);
nand NAND2_3290(N10928, N10873, 1'b1);
not NOT1_3314(N10988, N10928);
nand NAND2_3315(N10989, N10928, 1'b1);
nand NAND2_3350(N11044, N10989, 1'b1);
not NOT1_3380(N11114, N11044);
nand NAND2_3381(N11115, N11044, 1'b1);
nand NAND2_3410(N11168, N11115, 1'b1);
not NOT1_3425(N11213, N11168);
nand NAND2_3426(N11214, N11168, 1'b1);
nand NAND2_3446(N11242, N11213, 1'b1);
nand NAND2_3454(N11260, N11242, 1'b1);
and AND2_3466(N11278, N11260, 1'b1);
or OR2_3485(N11299, N11278, 1'b0);
nand NAND2_3491(N11313, N11299, 1'b1);
not NOT1_3492(N11314, N11299);
nand NAND2_3497(N11321, N11314, 1'b1);
nand NAND2_3500(N11328, N11321, 1'b1);
not NOT1_3504(N11334, N11328);

endmodule
