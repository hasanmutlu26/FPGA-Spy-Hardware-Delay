library verilog;
use verilog.vl_types.all;
entity delay_testbench is
end delay_testbench;
