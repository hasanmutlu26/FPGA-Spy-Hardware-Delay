library verilog;
use verilog.vl_types.all;
entity singlepath_plode_testbench is
end singlepath_plode_testbench;
