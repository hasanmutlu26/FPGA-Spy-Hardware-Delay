// Path to be chained: ro_18
// The path works as NOT: n
// Chain amount: 100

module ro_18_100(pathResult, pathInput);
input pathInput;
output pathResult;

(* keep = 1 *) wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98;

ro_18 p0(w0, pathInput);
ro_18 p1(w1, w0);
ro_18 p2(w2, w1);
ro_18 p3(w3, w2);
ro_18 p4(w4, w3);
ro_18 p5(w5, w4);
ro_18 p6(w6, w5);
ro_18 p7(w7, w6);
ro_18 p8(w8, w7);
ro_18 p9(w9, w8);
ro_18 p10(w10, w9);
ro_18 p11(w11, w10);
ro_18 p12(w12, w11);
ro_18 p13(w13, w12);
ro_18 p14(w14, w13);
ro_18 p15(w15, w14);
ro_18 p16(w16, w15);
ro_18 p17(w17, w16);
ro_18 p18(w18, w17);
ro_18 p19(w19, w18);
ro_18 p20(w20, w19);
ro_18 p21(w21, w20);
ro_18 p22(w22, w21);
ro_18 p23(w23, w22);
ro_18 p24(w24, w23);
ro_18 p25(w25, w24);
ro_18 p26(w26, w25);
ro_18 p27(w27, w26);
ro_18 p28(w28, w27);
ro_18 p29(w29, w28);
ro_18 p30(w30, w29);
ro_18 p31(w31, w30);
ro_18 p32(w32, w31);
ro_18 p33(w33, w32);
ro_18 p34(w34, w33);
ro_18 p35(w35, w34);
ro_18 p36(w36, w35);
ro_18 p37(w37, w36);
ro_18 p38(w38, w37);
ro_18 p39(w39, w38);
ro_18 p40(w40, w39);
ro_18 p41(w41, w40);
ro_18 p42(w42, w41);
ro_18 p43(w43, w42);
ro_18 p44(w44, w43);
ro_18 p45(w45, w44);
ro_18 p46(w46, w45);
ro_18 p47(w47, w46);
ro_18 p48(w48, w47);
ro_18 p49(w49, w48);
ro_18 p50(w50, w49);
ro_18 p51(w51, w50);
ro_18 p52(w52, w51);
ro_18 p53(w53, w52);
ro_18 p54(w54, w53);
ro_18 p55(w55, w54);
ro_18 p56(w56, w55);
ro_18 p57(w57, w56);
ro_18 p58(w58, w57);
ro_18 p59(w59, w58);
ro_18 p60(w60, w59);
ro_18 p61(w61, w60);
ro_18 p62(w62, w61);
ro_18 p63(w63, w62);
ro_18 p64(w64, w63);
ro_18 p65(w65, w64);
ro_18 p66(w66, w65);
ro_18 p67(w67, w66);
ro_18 p68(w68, w67);
ro_18 p69(w69, w68);
ro_18 p70(w70, w69);
ro_18 p71(w71, w70);
ro_18 p72(w72, w71);
ro_18 p73(w73, w72);
ro_18 p74(w74, w73);
ro_18 p75(w75, w74);
ro_18 p76(w76, w75);
ro_18 p77(w77, w76);
ro_18 p78(w78, w77);
ro_18 p79(w79, w78);
ro_18 p80(w80, w79);
ro_18 p81(w81, w80);
ro_18 p82(w82, w81);
ro_18 p83(w83, w82);
ro_18 p84(w84, w83);
ro_18 p85(w85, w84);
ro_18 p86(w86, w85);
ro_18 p87(w87, w86);
ro_18 p88(w88, w87);
ro_18 p89(w89, w88);
ro_18 p90(w90, w89);
ro_18 p91(w91, w90);
ro_18 p92(w92, w91);
ro_18 p93(w93, w92);
ro_18 p94(w94, w93);
ro_18 p95(w95, w94);
ro_18 p96(w96, w95);
ro_18 p97(w97, w96);
ro_18 p98(w98, w97);
ro_18 p99(pathResult, w98);

endmodule