library verilog;
use verilog.vl_types.all;
entity path1_testbench is
end path1_testbench;
