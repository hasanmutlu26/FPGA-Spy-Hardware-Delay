library verilog;
use verilog.vl_types.all;
entity path1 is
    port(
        \out\           : out    vl_logic;
        \in\            : in     vl_logic;
        w0              : out    vl_logic;
        w1              : out    vl_logic;
        w2              : out    vl_logic;
        w3              : out    vl_logic;
        w4              : out    vl_logic;
        w5              : out    vl_logic;
        w6              : out    vl_logic;
        w7              : out    vl_logic;
        w8              : out    vl_logic;
        w9              : out    vl_logic;
        w10             : out    vl_logic;
        w11             : out    vl_logic;
        w12             : out    vl_logic;
        w13             : out    vl_logic;
        w14             : out    vl_logic;
        w15             : out    vl_logic;
        w16             : out    vl_logic;
        w17             : out    vl_logic;
        w18             : out    vl_logic;
        w19             : out    vl_logic;
        w20             : out    vl_logic;
        w21             : out    vl_logic;
        w22             : out    vl_logic;
        w23             : out    vl_logic;
        w24             : out    vl_logic;
        w25             : out    vl_logic;
        w26             : out    vl_logic;
        w27             : out    vl_logic;
        w28             : out    vl_logic;
        w29             : out    vl_logic;
        w30             : out    vl_logic;
        w31             : out    vl_logic;
        w32             : out    vl_logic;
        w33             : out    vl_logic;
        w34             : out    vl_logic;
        w35             : out    vl_logic;
        w36             : out    vl_logic;
        w37             : out    vl_logic;
        w38             : out    vl_logic;
        w39             : out    vl_logic;
        w40             : out    vl_logic;
        w41             : out    vl_logic;
        w42             : out    vl_logic;
        w43             : out    vl_logic;
        w44             : out    vl_logic;
        w45             : out    vl_logic;
        w46             : out    vl_logic;
        w47             : out    vl_logic;
        w48             : out    vl_logic;
        w49             : out    vl_logic;
        w50             : out    vl_logic;
        w51             : out    vl_logic;
        w52             : out    vl_logic;
        w53             : out    vl_logic;
        w54             : out    vl_logic;
        w55             : out    vl_logic;
        w56             : out    vl_logic;
        w57             : out    vl_logic;
        w58             : out    vl_logic;
        w59             : out    vl_logic;
        w60             : out    vl_logic;
        w61             : out    vl_logic;
        w62             : out    vl_logic;
        w63             : out    vl_logic;
        w64             : out    vl_logic;
        w65             : out    vl_logic;
        w66             : out    vl_logic;
        w67             : out    vl_logic;
        w68             : out    vl_logic;
        w69             : out    vl_logic;
        w70             : out    vl_logic;
        w71             : out    vl_logic;
        w72             : out    vl_logic;
        w73             : out    vl_logic;
        w74             : out    vl_logic;
        w75             : out    vl_logic;
        w76             : out    vl_logic;
        w77             : out    vl_logic;
        w78             : out    vl_logic;
        w79             : out    vl_logic;
        w80             : out    vl_logic;
        w81             : out    vl_logic;
        w82             : out    vl_logic;
        w83             : out    vl_logic;
        w84             : out    vl_logic;
        w85             : out    vl_logic;
        w86             : out    vl_logic;
        w87             : out    vl_logic;
        w88             : out    vl_logic;
        w89             : out    vl_logic;
        w90             : out    vl_logic;
        w91             : out    vl_logic;
        w92             : out    vl_logic;
        w93             : out    vl_logic;
        w94             : out    vl_logic;
        w95             : out    vl_logic;
        w96             : out    vl_logic;
        w97             : out    vl_logic;
        w98             : out    vl_logic;
        w99             : out    vl_logic;
        w100            : out    vl_logic;
        w101            : out    vl_logic;
        w102            : out    vl_logic;
        w103            : out    vl_logic;
        w104            : out    vl_logic;
        w105            : out    vl_logic;
        w106            : out    vl_logic;
        w107            : out    vl_logic;
        w108            : out    vl_logic;
        w109            : out    vl_logic;
        w110            : out    vl_logic;
        w111            : out    vl_logic;
        w112            : out    vl_logic;
        w113            : out    vl_logic;
        w114            : out    vl_logic;
        w115            : out    vl_logic;
        w116            : out    vl_logic;
        w117            : out    vl_logic;
        w118            : out    vl_logic;
        w119            : out    vl_logic;
        w120            : out    vl_logic;
        w121            : out    vl_logic;
        w122            : out    vl_logic;
        w123            : out    vl_logic;
        w124            : out    vl_logic;
        w125            : out    vl_logic;
        w126            : out    vl_logic;
        w127            : out    vl_logic;
        w128            : out    vl_logic;
        w129            : out    vl_logic;
        w130            : out    vl_logic;
        w131            : out    vl_logic;
        w132            : out    vl_logic;
        w133            : out    vl_logic;
        w134            : out    vl_logic;
        w135            : out    vl_logic;
        w136            : out    vl_logic;
        w137            : out    vl_logic;
        w138            : out    vl_logic;
        w139            : out    vl_logic;
        w140            : out    vl_logic;
        w141            : out    vl_logic;
        w142            : out    vl_logic;
        w143            : out    vl_logic;
        w144            : out    vl_logic;
        w145            : out    vl_logic;
        w146            : out    vl_logic;
        w147            : out    vl_logic;
        w148            : out    vl_logic;
        w149            : out    vl_logic;
        w150            : out    vl_logic;
        w151            : out    vl_logic;
        w152            : out    vl_logic;
        w153            : out    vl_logic;
        w154            : out    vl_logic;
        w155            : out    vl_logic;
        w156            : out    vl_logic;
        w157            : out    vl_logic;
        w158            : out    vl_logic;
        w159            : out    vl_logic;
        w160            : out    vl_logic;
        w161            : out    vl_logic;
        w162            : out    vl_logic;
        w163            : out    vl_logic;
        w164            : out    vl_logic;
        w165            : out    vl_logic;
        w166            : out    vl_logic;
        w167            : out    vl_logic;
        w168            : out    vl_logic;
        w169            : out    vl_logic;
        w170            : out    vl_logic;
        w171            : out    vl_logic;
        w172            : out    vl_logic;
        w173            : out    vl_logic;
        w174            : out    vl_logic;
        w175            : out    vl_logic;
        w176            : out    vl_logic;
        w177            : out    vl_logic;
        w178            : out    vl_logic;
        w179            : out    vl_logic;
        w180            : out    vl_logic;
        w181            : out    vl_logic;
        w182            : out    vl_logic;
        w183            : out    vl_logic;
        w184            : out    vl_logic;
        w185            : out    vl_logic;
        w186            : out    vl_logic;
        w187            : out    vl_logic;
        w188            : out    vl_logic;
        w189            : out    vl_logic;
        w190            : out    vl_logic;
        w191            : out    vl_logic;
        w192            : out    vl_logic;
        w193            : out    vl_logic;
        w194            : out    vl_logic;
        w195            : out    vl_logic;
        w196            : out    vl_logic;
        w197            : out    vl_logic;
        w198            : out    vl_logic;
        w199            : out    vl_logic;
        w200            : out    vl_logic;
        w201            : out    vl_logic;
        w202            : out    vl_logic;
        w203            : out    vl_logic;
        w204            : out    vl_logic;
        w205            : out    vl_logic;
        w206            : out    vl_logic;
        w207            : out    vl_logic;
        w208            : out    vl_logic;
        w209            : out    vl_logic;
        w210            : out    vl_logic;
        w211            : out    vl_logic;
        w212            : out    vl_logic;
        w213            : out    vl_logic;
        w214            : out    vl_logic;
        w215            : out    vl_logic;
        w216            : out    vl_logic;
        w217            : out    vl_logic;
        w218            : out    vl_logic;
        w219            : out    vl_logic;
        w220            : out    vl_logic;
        w221            : out    vl_logic;
        w222            : out    vl_logic;
        w223            : out    vl_logic;
        w224            : out    vl_logic;
        w225            : out    vl_logic;
        w226            : out    vl_logic;
        w227            : out    vl_logic;
        w228            : out    vl_logic;
        w229            : out    vl_logic;
        w230            : out    vl_logic;
        w231            : out    vl_logic;
        w232            : out    vl_logic;
        w233            : out    vl_logic;
        w234            : out    vl_logic;
        w235            : out    vl_logic;
        w236            : out    vl_logic;
        w237            : out    vl_logic;
        w238            : out    vl_logic;
        w239            : out    vl_logic;
        w240            : out    vl_logic;
        w241            : out    vl_logic;
        w242            : out    vl_logic;
        w243            : out    vl_logic;
        w244            : out    vl_logic;
        w245            : out    vl_logic;
        w246            : out    vl_logic;
        w247            : out    vl_logic;
        w248            : out    vl_logic;
        w249            : out    vl_logic;
        w250            : out    vl_logic;
        w251            : out    vl_logic;
        w252            : out    vl_logic;
        w253            : out    vl_logic;
        w254            : out    vl_logic;
        w255            : out    vl_logic;
        w256            : out    vl_logic;
        w257            : out    vl_logic;
        w258            : out    vl_logic;
        w259            : out    vl_logic;
        w260            : out    vl_logic;
        w261            : out    vl_logic;
        w262            : out    vl_logic;
        w263            : out    vl_logic;
        w264            : out    vl_logic;
        w265            : out    vl_logic;
        w266            : out    vl_logic;
        w267            : out    vl_logic;
        w268            : out    vl_logic;
        w269            : out    vl_logic;
        w270            : out    vl_logic;
        w271            : out    vl_logic;
        w272            : out    vl_logic;
        w273            : out    vl_logic;
        w274            : out    vl_logic;
        w275            : out    vl_logic;
        w276            : out    vl_logic;
        w277            : out    vl_logic;
        w278            : out    vl_logic;
        w279            : out    vl_logic;
        w280            : out    vl_logic;
        w281            : out    vl_logic;
        w282            : out    vl_logic;
        w283            : out    vl_logic;
        w284            : out    vl_logic;
        w285            : out    vl_logic;
        w286            : out    vl_logic;
        w287            : out    vl_logic;
        w288            : out    vl_logic;
        w289            : out    vl_logic;
        w290            : out    vl_logic;
        w291            : out    vl_logic;
        w292            : out    vl_logic;
        w293            : out    vl_logic;
        w294            : out    vl_logic;
        w295            : out    vl_logic;
        w296            : out    vl_logic;
        w297            : out    vl_logic;
        w298            : out    vl_logic;
        w299            : out    vl_logic;
        w300            : out    vl_logic;
        w301            : out    vl_logic;
        w302            : out    vl_logic;
        w303            : out    vl_logic;
        w304            : out    vl_logic;
        w305            : out    vl_logic;
        w306            : out    vl_logic;
        w307            : out    vl_logic;
        w308            : out    vl_logic;
        w309            : out    vl_logic;
        w310            : out    vl_logic;
        w311            : out    vl_logic;
        w312            : out    vl_logic;
        w313            : out    vl_logic;
        w314            : out    vl_logic;
        w315            : out    vl_logic;
        w316            : out    vl_logic;
        w317            : out    vl_logic;
        w318            : out    vl_logic;
        w319            : out    vl_logic;
        w320            : out    vl_logic;
        w321            : out    vl_logic;
        w322            : out    vl_logic;
        w323            : out    vl_logic;
        w324            : out    vl_logic;
        w325            : out    vl_logic;
        w326            : out    vl_logic;
        w327            : out    vl_logic;
        w328            : out    vl_logic;
        w329            : out    vl_logic;
        w330            : out    vl_logic;
        w331            : out    vl_logic;
        w332            : out    vl_logic;
        w333            : out    vl_logic;
        w334            : out    vl_logic;
        w335            : out    vl_logic;
        w336            : out    vl_logic;
        w337            : out    vl_logic;
        w338            : out    vl_logic;
        w339            : out    vl_logic;
        w340            : out    vl_logic;
        w341            : out    vl_logic;
        w342            : out    vl_logic;
        w343            : out    vl_logic;
        w344            : out    vl_logic;
        w345            : out    vl_logic;
        w346            : out    vl_logic;
        w347            : out    vl_logic;
        w348            : out    vl_logic;
        w349            : out    vl_logic;
        w350            : out    vl_logic;
        w351            : out    vl_logic;
        w352            : out    vl_logic;
        w353            : out    vl_logic;
        w354            : out    vl_logic;
        w355            : out    vl_logic;
        w356            : out    vl_logic;
        w357            : out    vl_logic;
        w358            : out    vl_logic;
        w359            : out    vl_logic;
        w360            : out    vl_logic;
        w361            : out    vl_logic;
        w362            : out    vl_logic;
        w363            : out    vl_logic;
        w364            : out    vl_logic;
        w365            : out    vl_logic;
        w366            : out    vl_logic;
        w367            : out    vl_logic;
        w368            : out    vl_logic;
        w369            : out    vl_logic;
        w370            : out    vl_logic;
        w371            : out    vl_logic;
        w372            : out    vl_logic;
        w373            : out    vl_logic;
        w374            : out    vl_logic;
        w375            : out    vl_logic;
        w376            : out    vl_logic;
        w377            : out    vl_logic;
        w378            : out    vl_logic;
        w379            : out    vl_logic;
        w380            : out    vl_logic;
        w381            : out    vl_logic;
        w382            : out    vl_logic;
        w383            : out    vl_logic;
        w384            : out    vl_logic;
        w385            : out    vl_logic;
        w386            : out    vl_logic;
        w387            : out    vl_logic;
        w388            : out    vl_logic;
        w389            : out    vl_logic;
        w390            : out    vl_logic;
        w391            : out    vl_logic;
        w392            : out    vl_logic;
        w393            : out    vl_logic;
        w394            : out    vl_logic;
        w395            : out    vl_logic;
        w396            : out    vl_logic;
        w397            : out    vl_logic;
        w398            : out    vl_logic;
        w399            : out    vl_logic;
        w400            : out    vl_logic;
        w401            : out    vl_logic;
        w402            : out    vl_logic;
        w403            : out    vl_logic;
        w404            : out    vl_logic;
        w405            : out    vl_logic;
        w406            : out    vl_logic;
        w407            : out    vl_logic;
        w408            : out    vl_logic;
        w409            : out    vl_logic;
        w410            : out    vl_logic;
        w411            : out    vl_logic;
        w412            : out    vl_logic;
        w413            : out    vl_logic;
        w414            : out    vl_logic;
        w415            : out    vl_logic;
        w416            : out    vl_logic;
        w417            : out    vl_logic;
        w418            : out    vl_logic;
        w419            : out    vl_logic;
        w420            : out    vl_logic;
        w421            : out    vl_logic;
        w422            : out    vl_logic;
        w423            : out    vl_logic;
        w424            : out    vl_logic;
        w425            : out    vl_logic;
        w426            : out    vl_logic;
        w427            : out    vl_logic;
        w428            : out    vl_logic;
        w429            : out    vl_logic;
        w430            : out    vl_logic;
        w431            : out    vl_logic;
        w432            : out    vl_logic;
        w433            : out    vl_logic;
        w434            : out    vl_logic;
        w435            : out    vl_logic;
        w436            : out    vl_logic;
        w437            : out    vl_logic;
        w438            : out    vl_logic;
        w439            : out    vl_logic;
        w440            : out    vl_logic;
        w441            : out    vl_logic;
        w442            : out    vl_logic;
        w443            : out    vl_logic;
        w444            : out    vl_logic;
        w445            : out    vl_logic;
        w446            : out    vl_logic;
        w447            : out    vl_logic;
        w448            : out    vl_logic;
        w449            : out    vl_logic;
        w450            : out    vl_logic;
        w451            : out    vl_logic;
        w452            : out    vl_logic;
        w453            : out    vl_logic;
        w454            : out    vl_logic;
        w455            : out    vl_logic;
        w456            : out    vl_logic;
        w457            : out    vl_logic;
        w458            : out    vl_logic;
        w459            : out    vl_logic;
        w460            : out    vl_logic;
        w461            : out    vl_logic;
        w462            : out    vl_logic;
        w463            : out    vl_logic;
        w464            : out    vl_logic;
        w465            : out    vl_logic;
        w466            : out    vl_logic;
        w467            : out    vl_logic;
        w468            : out    vl_logic;
        w469            : out    vl_logic;
        w470            : out    vl_logic;
        w471            : out    vl_logic;
        w472            : out    vl_logic;
        w473            : out    vl_logic;
        w474            : out    vl_logic;
        w475            : out    vl_logic;
        w476            : out    vl_logic;
        w477            : out    vl_logic;
        w478            : out    vl_logic;
        w479            : out    vl_logic;
        w480            : out    vl_logic;
        w481            : out    vl_logic;
        w482            : out    vl_logic;
        w483            : out    vl_logic;
        w484            : out    vl_logic;
        w485            : out    vl_logic;
        w486            : out    vl_logic;
        w487            : out    vl_logic;
        w488            : out    vl_logic;
        w489            : out    vl_logic;
        w490            : out    vl_logic;
        w491            : out    vl_logic;
        w492            : out    vl_logic;
        w493            : out    vl_logic;
        w494            : out    vl_logic;
        w495            : out    vl_logic;
        w496            : out    vl_logic;
        w497            : out    vl_logic;
        w498            : out    vl_logic;
        w499            : out    vl_logic;
        w500            : out    vl_logic;
        w501            : out    vl_logic;
        w502            : out    vl_logic;
        w503            : out    vl_logic;
        w504            : out    vl_logic;
        w505            : out    vl_logic;
        w506            : out    vl_logic;
        w507            : out    vl_logic;
        w508            : out    vl_logic;
        w509            : out    vl_logic;
        w510            : out    vl_logic;
        w511            : out    vl_logic;
        w512            : out    vl_logic;
        w513            : out    vl_logic;
        w514            : out    vl_logic;
        w515            : out    vl_logic;
        w516            : out    vl_logic;
        w517            : out    vl_logic;
        w518            : out    vl_logic;
        w519            : out    vl_logic;
        w520            : out    vl_logic;
        w521            : out    vl_logic;
        w522            : out    vl_logic;
        w523            : out    vl_logic;
        w524            : out    vl_logic;
        w525            : out    vl_logic;
        w526            : out    vl_logic;
        w527            : out    vl_logic;
        w528            : out    vl_logic;
        w529            : out    vl_logic;
        w530            : out    vl_logic;
        w531            : out    vl_logic;
        w532            : out    vl_logic;
        w533            : out    vl_logic;
        w534            : out    vl_logic;
        w535            : out    vl_logic;
        w536            : out    vl_logic;
        w537            : out    vl_logic;
        w538            : out    vl_logic;
        w539            : out    vl_logic;
        w540            : out    vl_logic;
        w541            : out    vl_logic;
        w542            : out    vl_logic;
        w543            : out    vl_logic;
        w544            : out    vl_logic;
        w545            : out    vl_logic;
        w546            : out    vl_logic;
        w547            : out    vl_logic;
        w548            : out    vl_logic;
        w549            : out    vl_logic;
        w550            : out    vl_logic;
        w551            : out    vl_logic;
        w552            : out    vl_logic;
        w553            : out    vl_logic;
        w554            : out    vl_logic;
        w555            : out    vl_logic;
        w556            : out    vl_logic;
        w557            : out    vl_logic;
        w558            : out    vl_logic;
        w559            : out    vl_logic;
        w560            : out    vl_logic;
        w561            : out    vl_logic;
        w562            : out    vl_logic;
        w563            : out    vl_logic;
        w564            : out    vl_logic;
        w565            : out    vl_logic;
        w566            : out    vl_logic;
        w567            : out    vl_logic;
        w568            : out    vl_logic;
        w569            : out    vl_logic;
        w570            : out    vl_logic;
        w571            : out    vl_logic;
        w572            : out    vl_logic;
        w573            : out    vl_logic;
        w574            : out    vl_logic;
        w575            : out    vl_logic;
        w576            : out    vl_logic;
        w577            : out    vl_logic;
        w578            : out    vl_logic;
        w579            : out    vl_logic;
        w580            : out    vl_logic;
        w581            : out    vl_logic;
        w582            : out    vl_logic;
        w583            : out    vl_logic;
        w584            : out    vl_logic;
        w585            : out    vl_logic;
        w586            : out    vl_logic;
        w587            : out    vl_logic;
        w588            : out    vl_logic;
        w589            : out    vl_logic;
        w590            : out    vl_logic;
        w591            : out    vl_logic;
        w592            : out    vl_logic;
        w593            : out    vl_logic;
        w594            : out    vl_logic;
        w595            : out    vl_logic;
        w596            : out    vl_logic;
        w597            : out    vl_logic;
        w598            : out    vl_logic;
        w599            : out    vl_logic;
        w600            : out    vl_logic;
        w601            : out    vl_logic;
        w602            : out    vl_logic;
        w603            : out    vl_logic;
        w604            : out    vl_logic;
        w605            : out    vl_logic;
        w606            : out    vl_logic;
        w607            : out    vl_logic;
        w608            : out    vl_logic;
        w609            : out    vl_logic;
        w610            : out    vl_logic;
        w611            : out    vl_logic;
        w612            : out    vl_logic;
        w613            : out    vl_logic;
        w614            : out    vl_logic;
        w615            : out    vl_logic;
        w616            : out    vl_logic;
        w617            : out    vl_logic;
        w618            : out    vl_logic;
        w619            : out    vl_logic;
        w620            : out    vl_logic;
        w621            : out    vl_logic;
        w622            : out    vl_logic;
        w623            : out    vl_logic;
        w624            : out    vl_logic;
        w625            : out    vl_logic;
        w626            : out    vl_logic;
        w627            : out    vl_logic;
        w628            : out    vl_logic;
        w629            : out    vl_logic;
        w630            : out    vl_logic;
        w631            : out    vl_logic;
        w632            : out    vl_logic;
        w633            : out    vl_logic;
        w634            : out    vl_logic;
        w635            : out    vl_logic;
        w636            : out    vl_logic;
        w637            : out    vl_logic;
        w638            : out    vl_logic;
        w639            : out    vl_logic;
        w640            : out    vl_logic;
        w641            : out    vl_logic;
        w642            : out    vl_logic;
        w643            : out    vl_logic;
        w644            : out    vl_logic;
        w645            : out    vl_logic;
        w646            : out    vl_logic;
        w647            : out    vl_logic;
        w648            : out    vl_logic;
        w649            : out    vl_logic;
        w650            : out    vl_logic;
        w651            : out    vl_logic;
        w652            : out    vl_logic;
        w653            : out    vl_logic;
        w654            : out    vl_logic;
        w655            : out    vl_logic;
        w656            : out    vl_logic;
        w657            : out    vl_logic;
        w658            : out    vl_logic;
        w659            : out    vl_logic;
        w660            : out    vl_logic;
        w661            : out    vl_logic;
        w662            : out    vl_logic;
        w663            : out    vl_logic;
        w664            : out    vl_logic;
        w665            : out    vl_logic;
        w666            : out    vl_logic;
        w667            : out    vl_logic;
        w668            : out    vl_logic;
        w669            : out    vl_logic;
        w670            : out    vl_logic;
        w671            : out    vl_logic;
        w672            : out    vl_logic;
        w673            : out    vl_logic;
        w674            : out    vl_logic;
        w675            : out    vl_logic;
        w676            : out    vl_logic;
        w677            : out    vl_logic;
        w678            : out    vl_logic;
        w679            : out    vl_logic;
        w680            : out    vl_logic;
        w681            : out    vl_logic;
        w682            : out    vl_logic;
        w683            : out    vl_logic;
        w684            : out    vl_logic;
        w685            : out    vl_logic;
        w686            : out    vl_logic;
        w687            : out    vl_logic;
        w688            : out    vl_logic;
        w689            : out    vl_logic;
        w690            : out    vl_logic;
        w691            : out    vl_logic;
        w692            : out    vl_logic;
        w693            : out    vl_logic;
        w694            : out    vl_logic;
        w695            : out    vl_logic;
        w696            : out    vl_logic;
        w697            : out    vl_logic;
        w698            : out    vl_logic;
        w699            : out    vl_logic;
        w700            : out    vl_logic;
        w701            : out    vl_logic;
        w702            : out    vl_logic;
        w703            : out    vl_logic;
        w704            : out    vl_logic;
        w705            : out    vl_logic;
        w706            : out    vl_logic;
        w707            : out    vl_logic;
        w708            : out    vl_logic;
        w709            : out    vl_logic;
        w710            : out    vl_logic;
        w711            : out    vl_logic;
        w712            : out    vl_logic;
        w713            : out    vl_logic;
        w714            : out    vl_logic;
        w715            : out    vl_logic;
        w716            : out    vl_logic;
        w717            : out    vl_logic;
        w718            : out    vl_logic;
        w719            : out    vl_logic;
        w720            : out    vl_logic;
        w721            : out    vl_logic;
        w722            : out    vl_logic;
        w723            : out    vl_logic;
        w724            : out    vl_logic;
        w725            : out    vl_logic;
        w726            : out    vl_logic;
        w727            : out    vl_logic;
        w728            : out    vl_logic;
        w729            : out    vl_logic;
        w730            : out    vl_logic;
        w731            : out    vl_logic;
        w732            : out    vl_logic;
        w733            : out    vl_logic;
        w734            : out    vl_logic;
        w735            : out    vl_logic;
        w736            : out    vl_logic;
        w737            : out    vl_logic;
        w738            : out    vl_logic;
        w739            : out    vl_logic;
        w740            : out    vl_logic;
        w741            : out    vl_logic;
        w742            : out    vl_logic;
        w743            : out    vl_logic;
        w744            : out    vl_logic;
        w745            : out    vl_logic;
        w746            : out    vl_logic;
        w747            : out    vl_logic;
        w748            : out    vl_logic;
        w749            : out    vl_logic;
        w750            : out    vl_logic;
        w751            : out    vl_logic;
        w752            : out    vl_logic;
        w753            : out    vl_logic;
        w754            : out    vl_logic;
        w755            : out    vl_logic;
        w756            : out    vl_logic;
        w757            : out    vl_logic;
        w758            : out    vl_logic;
        w759            : out    vl_logic;
        w760            : out    vl_logic;
        w761            : out    vl_logic;
        w762            : out    vl_logic;
        w763            : out    vl_logic;
        w764            : out    vl_logic;
        w765            : out    vl_logic;
        w766            : out    vl_logic;
        w767            : out    vl_logic;
        w768            : out    vl_logic;
        w769            : out    vl_logic;
        w770            : out    vl_logic;
        w771            : out    vl_logic;
        w772            : out    vl_logic;
        w773            : out    vl_logic;
        w774            : out    vl_logic;
        w775            : out    vl_logic;
        w776            : out    vl_logic;
        w777            : out    vl_logic;
        w778            : out    vl_logic;
        w779            : out    vl_logic;
        w780            : out    vl_logic;
        w781            : out    vl_logic;
        w782            : out    vl_logic;
        w783            : out    vl_logic;
        w784            : out    vl_logic;
        w785            : out    vl_logic;
        w786            : out    vl_logic;
        w787            : out    vl_logic;
        w788            : out    vl_logic;
        w789            : out    vl_logic;
        w790            : out    vl_logic;
        w791            : out    vl_logic;
        w792            : out    vl_logic;
        w793            : out    vl_logic;
        w794            : out    vl_logic;
        w795            : out    vl_logic;
        w796            : out    vl_logic;
        w797            : out    vl_logic;
        w798            : out    vl_logic;
        w799            : out    vl_logic;
        w800            : out    vl_logic;
        w801            : out    vl_logic;
        w802            : out    vl_logic;
        w803            : out    vl_logic;
        w804            : out    vl_logic;
        w805            : out    vl_logic;
        w806            : out    vl_logic;
        w807            : out    vl_logic;
        w808            : out    vl_logic;
        w809            : out    vl_logic;
        w810            : out    vl_logic;
        w811            : out    vl_logic;
        w812            : out    vl_logic;
        w813            : out    vl_logic;
        w814            : out    vl_logic;
        w815            : out    vl_logic;
        w816            : out    vl_logic;
        w817            : out    vl_logic;
        w818            : out    vl_logic;
        w819            : out    vl_logic;
        w820            : out    vl_logic;
        w821            : out    vl_logic;
        w822            : out    vl_logic;
        w823            : out    vl_logic;
        w824            : out    vl_logic;
        w825            : out    vl_logic;
        w826            : out    vl_logic;
        w827            : out    vl_logic;
        w828            : out    vl_logic;
        w829            : out    vl_logic;
        w830            : out    vl_logic;
        w831            : out    vl_logic;
        w832            : out    vl_logic;
        w833            : out    vl_logic;
        w834            : out    vl_logic;
        w835            : out    vl_logic;
        w836            : out    vl_logic;
        w837            : out    vl_logic;
        w838            : out    vl_logic;
        w839            : out    vl_logic;
        w840            : out    vl_logic;
        w841            : out    vl_logic;
        w842            : out    vl_logic;
        w843            : out    vl_logic;
        w844            : out    vl_logic;
        w845            : out    vl_logic;
        w846            : out    vl_logic;
        w847            : out    vl_logic;
        w848            : out    vl_logic;
        w849            : out    vl_logic;
        w850            : out    vl_logic;
        w851            : out    vl_logic;
        w852            : out    vl_logic;
        w853            : out    vl_logic;
        w854            : out    vl_logic;
        w855            : out    vl_logic;
        w856            : out    vl_logic;
        w857            : out    vl_logic;
        w858            : out    vl_logic;
        w859            : out    vl_logic;
        w860            : out    vl_logic;
        w861            : out    vl_logic;
        w862            : out    vl_logic;
        w863            : out    vl_logic;
        w864            : out    vl_logic;
        w865            : out    vl_logic;
        w866            : out    vl_logic;
        w867            : out    vl_logic;
        w868            : out    vl_logic;
        w869            : out    vl_logic;
        w870            : out    vl_logic;
        w871            : out    vl_logic;
        w872            : out    vl_logic;
        w873            : out    vl_logic;
        w874            : out    vl_logic;
        w875            : out    vl_logic;
        w876            : out    vl_logic;
        w877            : out    vl_logic;
        w878            : out    vl_logic;
        w879            : out    vl_logic;
        w880            : out    vl_logic;
        w881            : out    vl_logic;
        w882            : out    vl_logic;
        w883            : out    vl_logic;
        w884            : out    vl_logic;
        w885            : out    vl_logic;
        w886            : out    vl_logic;
        w887            : out    vl_logic;
        w888            : out    vl_logic;
        w889            : out    vl_logic;
        w890            : out    vl_logic;
        w891            : out    vl_logic;
        w892            : out    vl_logic;
        w893            : out    vl_logic;
        w894            : out    vl_logic;
        w895            : out    vl_logic;
        w896            : out    vl_logic;
        w897            : out    vl_logic;
        w898            : out    vl_logic;
        w899            : out    vl_logic;
        w900            : out    vl_logic;
        w901            : out    vl_logic;
        w902            : out    vl_logic;
        w903            : out    vl_logic;
        w904            : out    vl_logic;
        w905            : out    vl_logic;
        w906            : out    vl_logic;
        w907            : out    vl_logic;
        w908            : out    vl_logic;
        w909            : out    vl_logic;
        w910            : out    vl_logic;
        w911            : out    vl_logic;
        w912            : out    vl_logic;
        w913            : out    vl_logic;
        w914            : out    vl_logic;
        w915            : out    vl_logic;
        w916            : out    vl_logic;
        w917            : out    vl_logic;
        w918            : out    vl_logic;
        w919            : out    vl_logic;
        w920            : out    vl_logic;
        w921            : out    vl_logic;
        w922            : out    vl_logic;
        w923            : out    vl_logic;
        w924            : out    vl_logic;
        w925            : out    vl_logic;
        w926            : out    vl_logic;
        w927            : out    vl_logic;
        w928            : out    vl_logic;
        w929            : out    vl_logic;
        w930            : out    vl_logic;
        w931            : out    vl_logic;
        w932            : out    vl_logic;
        w933            : out    vl_logic;
        w934            : out    vl_logic;
        w935            : out    vl_logic;
        w936            : out    vl_logic;
        w937            : out    vl_logic;
        w938            : out    vl_logic;
        w939            : out    vl_logic;
        w940            : out    vl_logic;
        w941            : out    vl_logic;
        w942            : out    vl_logic;
        w943            : out    vl_logic;
        w944            : out    vl_logic;
        w945            : out    vl_logic;
        w946            : out    vl_logic;
        w947            : out    vl_logic;
        w948            : out    vl_logic;
        w949            : out    vl_logic;
        w950            : out    vl_logic;
        w951            : out    vl_logic;
        w952            : out    vl_logic;
        w953            : out    vl_logic;
        w954            : out    vl_logic;
        w955            : out    vl_logic;
        w956            : out    vl_logic;
        w957            : out    vl_logic;
        w958            : out    vl_logic;
        w959            : out    vl_logic;
        w960            : out    vl_logic;
        w961            : out    vl_logic;
        w962            : out    vl_logic;
        w963            : out    vl_logic;
        w964            : out    vl_logic;
        w965            : out    vl_logic;
        w966            : out    vl_logic;
        w967            : out    vl_logic;
        w968            : out    vl_logic;
        w969            : out    vl_logic;
        w970            : out    vl_logic;
        w971            : out    vl_logic;
        w972            : out    vl_logic;
        w973            : out    vl_logic;
        w974            : out    vl_logic;
        w975            : out    vl_logic;
        w976            : out    vl_logic;
        w977            : out    vl_logic;
        w978            : out    vl_logic;
        w979            : out    vl_logic;
        w980            : out    vl_logic;
        w981            : out    vl_logic;
        w982            : out    vl_logic;
        w983            : out    vl_logic;
        w984            : out    vl_logic;
        w985            : out    vl_logic;
        w986            : out    vl_logic;
        w987            : out    vl_logic;
        w988            : out    vl_logic;
        w989            : out    vl_logic;
        w990            : out    vl_logic;
        w991            : out    vl_logic;
        w992            : out    vl_logic;
        w993            : out    vl_logic;
        w994            : out    vl_logic;
        w995            : out    vl_logic;
        w996            : out    vl_logic;
        w997            : out    vl_logic;
        w998            : out    vl_logic
    );
end path1;
