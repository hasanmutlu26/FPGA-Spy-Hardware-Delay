module not3_34_50(pathResult, pathInput);
input pathInput;
output pathResult;

(* keep = 1 *) wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49;

not3_34 p0(w0, pathInput);
not3_34 p1(w1, w0);
not3_34 p2(w2, w1);
not3_34 p3(w3, w2);
not3_34 p4(w4, w3);
not3_34 p5(w5, w4);
not3_34 p6(w6, w5);
not3_34 p7(w7, w6);
not3_34 p8(w8, w7);
not3_34 p9(w9, w8);
not3_34 p10(w10, w9);
not3_34 p11(w11, w10);
not3_34 p12(w12, w11);
not3_34 p13(w13, w12);
not3_34 p14(w14, w13);
not3_34 p15(w15, w14);
not3_34 p16(w16, w15);
not3_34 p17(w17, w16);
not3_34 p18(w18, w17);
not3_34 p19(w19, w18);
not3_34 p20(w20, w19);
not3_34 p21(w21, w20);
not3_34 p22(w22, w21);
not3_34 p23(w23, w22);
not3_34 p24(w24, w23);
not3_34 p25(w25, w24);
not3_34 p26(w26, w25);
not3_34 p27(w27, w26);
not3_34 p28(w28, w27);
not3_34 p29(w29, w28);
not3_34 p30(w30, w29);
not3_34 p31(w31, w30);
not3_34 p32(w32, w31);
not3_34 p33(w33, w32);
not3_34 p34(w34, w33);
not3_34 p35(w35, w34);
not3_34 p36(w36, w35);
not3_34 p37(w37, w36);
not3_34 p38(w38, w37);
not3_34 p39(w39, w38);
not3_34 p40(w40, w39);
not3_34 p41(w41, w40);
not3_34 p42(w42, w41);
not3_34 p43(w43, w42);
not3_34 p44(w44, w43);
not3_34 p45(w45, w44);
not3_34 p46(w46, w45);
not3_34 p47(w47, w46);
not3_34 p48(w48, w47);
not3_34 p49(pathResult, w48);

endmodule
