module singlepath_1_6.v(pathResult, pathInput);
input pathInput;
output pathResult;
(* keep = 1 *) wire 