library verilog;
use verilog.vl_types.all;
entity path2 is
    port(
        \out\           : out    vl_logic;
        \in\            : in     vl_logic
    );
end path2;
