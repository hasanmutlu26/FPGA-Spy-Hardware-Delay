module singlepath_3_wrapper(pathResult, pathInput);
(* keep = 1 *) input pathInput;
(* keep = 1 *) output pathResult;

(* keep = 1 *) wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98;

singlepath_3 p0(w0, pathInput);
singlepath_3 p1(w1, w0);
singlepath_3 p2(w2, w1);
singlepath_3 p3(w3, w2);
singlepath_3 p4(w4, w3);
singlepath_3 p5(w5, w4);
singlepath_3 p6(w6, w5);
singlepath_3 p7(w7, w6);
singlepath_3 p8(w8, w7);
singlepath_3 p9(w9, w8);
singlepath_3 p10(w10, w9);
singlepath_3 p11(w11, w10);
singlepath_3 p12(w12, w11);
singlepath_3 p13(w13, w12);
singlepath_3 p14(w14, w13);
singlepath_3 p15(w15, w14);
singlepath_3 p16(w16, w15);
singlepath_3 p17(w17, w16);
singlepath_3 p18(w18, w17);
singlepath_3 p19(w19, w18);
singlepath_3 p20(w20, w19);
singlepath_3 p21(w21, w20);
singlepath_3 p22(w22, w21);
singlepath_3 p23(w23, w22);
singlepath_3 p24(w24, w23);
singlepath_3 p25(w25, w24);
singlepath_3 p26(w26, w25);
singlepath_3 p27(w27, w26);
singlepath_3 p28(w28, w27);
singlepath_3 p29(w29, w28);
singlepath_3 p30(w30, w29);
singlepath_3 p31(w31, w30);
singlepath_3 p32(w32, w31);
singlepath_3 p33(w33, w32);
singlepath_3 p34(w34, w33);
singlepath_3 p35(w35, w34);
singlepath_3 p36(w36, w35);
singlepath_3 p37(w37, w36);
singlepath_3 p38(w38, w37);
singlepath_3 p39(w39, w38);
singlepath_3 p40(w40, w39);
singlepath_3 p41(w41, w40);
singlepath_3 p42(w42, w41);
singlepath_3 p43(w43, w42);
singlepath_3 p44(w44, w43);
singlepath_3 p45(w45, w44);
singlepath_3 p46(w46, w45);
singlepath_3 p47(w47, w46);
singlepath_3 p48(w48, w47);
singlepath_3 p49(pathResult, w48);
/*singlepath_3 p50(w50, w49);
singlepath_3 p51(w51, w50);
singlepath_3 p52(w52, w51);
singlepath_3 p53(w53, w52);
singlepath_3 p54(w54, w53);
singlepath_3 p55(w55, w54);
singlepath_3 p56(w56, w55);
singlepath_3 p57(w57, w56);
singlepath_3 p58(w58, w57);
singlepath_3 p59(w59, w58);
singlepath_3 p60(w60, w59);
singlepath_3 p61(w61, w60);
singlepath_3 p62(w62, w61);
singlepath_3 p63(w63, w62);
singlepath_3 p64(w64, w63);
singlepath_3 p65(w65, w64);
singlepath_3 p66(w66, w65);
singlepath_3 p67(w67, w66);
singlepath_3 p68(w68, w67);
singlepath_3 p69(w69, w68);
singlepath_3 p70(w70, w69);
singlepath_3 p71(w71, w70);
singlepath_3 p72(w72, w71);
singlepath_3 p73(w73, w72);
singlepath_3 p74(w74, w73);
singlepath_3 p75(w75, w74);
singlepath_3 p76(w76, w75);
singlepath_3 p77(w77, w76);
singlepath_3 p78(w78, w77);
singlepath_3 p79(w79, w78);
singlepath_3 p80(w80, w79);
singlepath_3 p81(w81, w80);
singlepath_3 p82(w82, w81);
singlepath_3 p83(w83, w82);
singlepath_3 p84(w84, w83);
singlepath_3 p85(w85, w84);
singlepath_3 p86(w86, w85);
singlepath_3 p87(w87, w86);
singlepath_3 p88(w88, w87);
singlepath_3 p89(w89, w88);
singlepath_3 p90(w90, w89);
singlepath_3 p91(w91, w90);
singlepath_3 p92(w92, w91);
singlepath_3 p93(w93, w92);
singlepath_3 p94(w94, w93);
singlepath_3 p95(w95, w94);
singlepath_3 p96(w96, w95);
singlepath_3 p97(w97, w96);
singlepath_3 p98(w98, w97);
singlepath_3 p99(pathResult, w98);*/


endmodule