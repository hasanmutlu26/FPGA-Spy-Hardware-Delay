
module not3_34_100(pathResult, pathInput);
input pathInput;
output pathResult;

(* keep = 1 *) wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98;
not3_34 p0(w0, pathInput);
not3_34 p1(w1, w0);
not3_34 p2(w2, w1);
not3_34 p3(w3, w2);
not3_34 p4(w4, w3);
not3_34 p5(w5, w4);
not3_34 p6(w6, w5);
not3_34 p7(w7, w6);
not3_34 p8(w8, w7);
not3_34 p9(w9, w8);
not3_34 p10(w10, w9);
not3_34 p11(w11, w10);
not3_34 p12(w12, w11);
not3_34 p13(w13, w12);
not3_34 p14(w14, w13);
not3_34 p15(w15, w14);
not3_34 p16(w16, w15);
not3_34 p17(w17, w16);
not3_34 p18(w18, w17);
not3_34 p19(w19, w18);
not3_34 p20(w20, w19);
not3_34 p21(w21, w20);
not3_34 p22(w22, w21);
not3_34 p23(w23, w22);
not3_34 p24(w24, w23);
not3_34 p25(w25, w24);
not3_34 p26(w26, w25);
not3_34 p27(w27, w26);
not3_34 p28(w28, w27);
not3_34 p29(w29, w28);
not3_34 p30(w30, w29);
not3_34 p31(w31, w30);
not3_34 p32(w32, w31);
not3_34 p33(w33, w32);
not3_34 p34(w34, w33);
not3_34 p35(w35, w34);
not3_34 p36(w36, w35);
not3_34 p37(w37, w36);
not3_34 p38(w38, w37);
not3_34 p39(w39, w38);
not3_34 p40(w40, w39);
not3_34 p41(w41, w40);
not3_34 p42(w42, w41);
not3_34 p43(w43, w42);
not3_34 p44(w44, w43);
not3_34 p45(w45, w44);
not3_34 p46(w46, w45);
not3_34 p47(w47, w46);
not3_34 p48(w48, w47);
not3_34 p49(w49, w48);
not3_34 p50(w50, w49);
not3_34 p51(w51, w50);
not3_34 p52(w52, w51);
not3_34 p53(w53, w52);
not3_34 p54(w54, w53);
not3_34 p55(w55, w54);
not3_34 p56(w56, w55);
not3_34 p57(w57, w56);
not3_34 p58(w58, w57);
not3_34 p59(w59, w58);
not3_34 p60(w60, w59);
not3_34 p61(w61, w60);
not3_34 p62(w62, w61);
not3_34 p63(w63, w62);
not3_34 p64(w64, w63);
not3_34 p65(w65, w64);
not3_34 p66(w66, w65);
not3_34 p67(w67, w66);
not3_34 p68(w68, w67);
not3_34 p69(w69, w68);
not3_34 p70(w70, w69);
not3_34 p71(w71, w70);
not3_34 p72(w72, w71);
not3_34 p73(w73, w72);
not3_34 p74(w74, w73);
not3_34 p75(w75, w74);
not3_34 p76(w76, w75);
not3_34 p77(w77, w76);
not3_34 p78(w78, w77);
not3_34 p79(w79, w78);
not3_34 p80(w80, w79);
not3_34 p81(w81, w80);
not3_34 p82(w82, w81);
not3_34 p83(w83, w82);
not3_34 p84(w84, w83);
not3_34 p85(w85, w84);
not3_34 p86(w86, w85);
not3_34 p87(w87, w86);
not3_34 p88(w88, w87);
not3_34 p89(w89, w88);
not3_34 p90(w90, w89);
not3_34 p91(w91, w90);
not3_34 p92(w92, w91);
not3_34 p93(w93, w92);
not3_34 p94(w94, w93);
not3_34 p95(w95, w94);
not3_34 p96(w96, w95);
not3_34 p97(w97, w96);
not3_34 p98(w98, w97);
not3_34 p99(pathResult, w98);

endmodule



