library verilog;
use verilog.vl_types.all;
entity singlepath_plode is
    port(
        N8076           : out    vl_logic;
        N411            : in     vl_logic;
        VCC             : in     vl_logic;
        GND             : in     vl_logic;
        s1              : out    vl_logic;
        s2              : out    vl_logic;
        s3              : out    vl_logic;
        s4              : out    vl_logic;
        s5              : out    vl_logic;
        s6              : out    vl_logic;
        s7              : out    vl_logic;
        s8              : out    vl_logic;
        s9              : out    vl_logic;
        s10             : out    vl_logic;
        s11             : out    vl_logic;
        s12             : out    vl_logic;
        s13             : out    vl_logic;
        s14             : out    vl_logic;
        s15             : out    vl_logic;
        s16             : out    vl_logic;
        s17             : out    vl_logic;
        s18             : out    vl_logic;
        s19             : out    vl_logic;
        s20             : out    vl_logic;
        s21             : out    vl_logic;
        s22             : out    vl_logic;
        s23             : out    vl_logic;
        s24             : out    vl_logic;
        s25             : out    vl_logic;
        s26             : out    vl_logic;
        s27             : out    vl_logic;
        s28             : out    vl_logic;
        s29             : out    vl_logic
    );
end singlepath_plode;
