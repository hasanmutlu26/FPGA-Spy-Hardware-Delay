// Path to be chained: ro_35n
// The path works as NOT: y
// Chain amount: 100

module ro_35n_100(pathResult, pathInput);
input pathInput;
output pathResult;

(* keep = 1 *) wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98;

ro_35n p0(w0, pathInput);
ro_35n p1(w1, w0);
ro_35n p2(w2, w1);
ro_35n p3(w3, w2);
ro_35n p4(w4, w3);
ro_35n p5(w5, w4);
ro_35n p6(w6, w5);
ro_35n p7(w7, w6);
ro_35n p8(w8, w7);
ro_35n p9(w9, w8);
ro_35n p10(w10, w9);
ro_35n p11(w11, w10);
ro_35n p12(w12, w11);
ro_35n p13(w13, w12);
ro_35n p14(w14, w13);
ro_35n p15(w15, w14);
ro_35n p16(w16, w15);
ro_35n p17(w17, w16);
ro_35n p18(w18, w17);
ro_35n p19(w19, w18);
ro_35n p20(w20, w19);
ro_35n p21(w21, w20);
ro_35n p22(w22, w21);
ro_35n p23(w23, w22);
ro_35n p24(w24, w23);
ro_35n p25(w25, w24);
ro_35n p26(w26, w25);
ro_35n p27(w27, w26);
ro_35n p28(w28, w27);
ro_35n p29(w29, w28);
ro_35n p30(w30, w29);
ro_35n p31(w31, w30);
ro_35n p32(w32, w31);
ro_35n p33(w33, w32);
ro_35n p34(w34, w33);
ro_35n p35(w35, w34);
ro_35n p36(w36, w35);
ro_35n p37(w37, w36);
ro_35n p38(w38, w37);
ro_35n p39(w39, w38);
ro_35n p40(w40, w39);
ro_35n p41(w41, w40);
ro_35n p42(w42, w41);
ro_35n p43(w43, w42);
ro_35n p44(w44, w43);
ro_35n p45(w45, w44);
ro_35n p46(w46, w45);
ro_35n p47(w47, w46);
ro_35n p48(w48, w47);
ro_35n p49(w49, w48);
ro_35n p50(w50, w49);
ro_35n p51(w51, w50);
ro_35n p52(w52, w51);
ro_35n p53(w53, w52);
ro_35n p54(w54, w53);
ro_35n p55(w55, w54);
ro_35n p56(w56, w55);
ro_35n p57(w57, w56);
ro_35n p58(w58, w57);
ro_35n p59(w59, w58);
ro_35n p60(w60, w59);
ro_35n p61(w61, w60);
ro_35n p62(w62, w61);
ro_35n p63(w63, w62);
ro_35n p64(w64, w63);
ro_35n p65(w65, w64);
ro_35n p66(w66, w65);
ro_35n p67(w67, w66);
ro_35n p68(w68, w67);
ro_35n p69(w69, w68);
ro_35n p70(w70, w69);
ro_35n p71(w71, w70);
ro_35n p72(w72, w71);
ro_35n p73(w73, w72);
ro_35n p74(w74, w73);
ro_35n p75(w75, w74);
ro_35n p76(w76, w75);
ro_35n p77(w77, w76);
ro_35n p78(w78, w77);
ro_35n p79(w79, w78);
ro_35n p80(w80, w79);
ro_35n p81(w81, w80);
ro_35n p82(w82, w81);
ro_35n p83(w83, w82);
ro_35n p84(w84, w83);
ro_35n p85(w85, w84);
ro_35n p86(w86, w85);
ro_35n p87(w87, w86);
ro_35n p88(w88, w87);
ro_35n p89(w89, w88);
ro_35n p90(w90, w89);
ro_35n p91(w91, w90);
ro_35n p92(w92, w91);
ro_35n p93(w93, w92);
ro_35n p94(w94, w93);
ro_35n p95(w95, w94);
ro_35n p96(w96, w95);
ro_35n p97(w97, w96);
ro_35n p98(w98, w97);
ro_35n p99(pathResult, w98);

endmodule