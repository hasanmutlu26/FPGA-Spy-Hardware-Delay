library verilog;
use verilog.vl_types.all;
entity HightoLow_testbench is
end HightoLow_testbench;
