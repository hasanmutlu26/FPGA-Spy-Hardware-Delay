// Path to be chained: ro_17n
// The path works as NOT: y
// Chain amount: 100

module ro_17n_100(pathResult, pathInput);
input pathInput;
output pathResult;

(* keep = 1 *) wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98;

ro_17n p0(w0, pathInput);
ro_17n p1(w1, w0);
ro_17n p2(w2, w1);
ro_17n p3(w3, w2);
ro_17n p4(w4, w3);
ro_17n p5(w5, w4);
ro_17n p6(w6, w5);
ro_17n p7(w7, w6);
ro_17n p8(w8, w7);
ro_17n p9(w9, w8);
ro_17n p10(w10, w9);
ro_17n p11(w11, w10);
ro_17n p12(w12, w11);
ro_17n p13(w13, w12);
ro_17n p14(w14, w13);
ro_17n p15(w15, w14);
ro_17n p16(w16, w15);
ro_17n p17(w17, w16);
ro_17n p18(w18, w17);
ro_17n p19(w19, w18);
ro_17n p20(w20, w19);
ro_17n p21(w21, w20);
ro_17n p22(w22, w21);
ro_17n p23(w23, w22);
ro_17n p24(w24, w23);
ro_17n p25(w25, w24);
ro_17n p26(w26, w25);
ro_17n p27(w27, w26);
ro_17n p28(w28, w27);
ro_17n p29(w29, w28);
ro_17n p30(w30, w29);
ro_17n p31(w31, w30);
ro_17n p32(w32, w31);
ro_17n p33(w33, w32);
ro_17n p34(w34, w33);
ro_17n p35(w35, w34);
ro_17n p36(w36, w35);
ro_17n p37(w37, w36);
ro_17n p38(w38, w37);
ro_17n p39(w39, w38);
ro_17n p40(w40, w39);
ro_17n p41(w41, w40);
ro_17n p42(w42, w41);
ro_17n p43(w43, w42);
ro_17n p44(w44, w43);
ro_17n p45(w45, w44);
ro_17n p46(w46, w45);
ro_17n p47(w47, w46);
ro_17n p48(w48, w47);
ro_17n p49(w49, w48);
ro_17n p50(w50, w49);
ro_17n p51(w51, w50);
ro_17n p52(w52, w51);
ro_17n p53(w53, w52);
ro_17n p54(w54, w53);
ro_17n p55(w55, w54);
ro_17n p56(w56, w55);
ro_17n p57(w57, w56);
ro_17n p58(w58, w57);
ro_17n p59(w59, w58);
ro_17n p60(w60, w59);
ro_17n p61(w61, w60);
ro_17n p62(w62, w61);
ro_17n p63(w63, w62);
ro_17n p64(w64, w63);
ro_17n p65(w65, w64);
ro_17n p66(w66, w65);
ro_17n p67(w67, w66);
ro_17n p68(w68, w67);
ro_17n p69(w69, w68);
ro_17n p70(w70, w69);
ro_17n p71(w71, w70);
ro_17n p72(w72, w71);
ro_17n p73(w73, w72);
ro_17n p74(w74, w73);
ro_17n p75(w75, w74);
ro_17n p76(w76, w75);
ro_17n p77(w77, w76);
ro_17n p78(w78, w77);
ro_17n p79(w79, w78);
ro_17n p80(w80, w79);
ro_17n p81(w81, w80);
ro_17n p82(w82, w81);
ro_17n p83(w83, w82);
ro_17n p84(w84, w83);
ro_17n p85(w85, w84);
ro_17n p86(w86, w85);
ro_17n p87(w87, w86);
ro_17n p88(w88, w87);
ro_17n p89(w89, w88);
ro_17n p90(w90, w89);
ro_17n p91(w91, w90);
ro_17n p92(w92, w91);
ro_17n p93(w93, w92);
ro_17n p94(w94, w93);
ro_17n p95(w95, w94);
ro_17n p96(w96, w95);
ro_17n p97(w97, w96);
ro_17n p98(w98, w97);
ro_17n p99(pathResult, w98);

endmodule