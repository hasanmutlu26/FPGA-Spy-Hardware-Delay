library verilog;
use verilog.vl_types.all;
entity decToSeg_testbench is
end decToSeg_testbench;
